parameter int COEFF_WIDTH = 16;
parameter int N_TAPS = 150;
parameter logic signed[COEFF_WIDTH-1:0] filter_coeffs[0:N_TAPS-1] = {
    16'b1111111111111001,
    16'b1111111111101110,
    16'b1111111111011101,
    16'b1111111111001000,
    16'b1111111110110111,
    16'b1111111110110011,
    16'b1111111111000110,
    16'b1111111111111000,
    16'b0000000001001101,
    16'b0000000010111011,
    16'b0000000100110010,
    16'b0000000110011000,
    16'b0000000111010010,
    16'b0000000111001110,
    16'b0000000110000110,
    16'b0000000100000101,
    16'b0000000001101001,
    16'b1111111111011000,
    16'b1111111101110111,
    16'b1111111101011101,
    16'b1111111110001101,
    16'b1111111111110000,
    16'b0000000001011111,
    16'b0000000010101111,
    16'b0000000011000010,
    16'b0000000010001110,
    16'b0000000000100110,
    16'b1111111110110000,
    16'b1111111101011010,
    16'b1111111101000111,
    16'b1111111110000000,
    16'b1111111111110001,
    16'b0000000001101110,
    16'b0000000011000100,
    16'b0000000011001101,
    16'b0000000010000001,
    16'b1111111111111011,
    16'b1111111101101111,
    16'b1111111100010111,
    16'b1111111100011100,
    16'b1111111110000010,
    16'b0000000000100101,
    16'b0000000011000101,
    16'b0000000100011101,
    16'b0000000100000011,
    16'b0000000001111001,
    16'b1111111110101110,
    16'b1111111011110101,
    16'b1111111010011110,
    16'b1111111011010110,
    16'b1111111110010101,
    16'b0000000010010100,
    16'b0000000101101110,
    16'b0000000111000001,
    16'b0000000101011010,
    16'b0000000001010001,
    16'b1111111100000100,
    16'b1111110111111011,
    16'b1111110110110010,
    16'b1111111001100010,
    16'b1111111111100100,
    16'b0000000110101111,
    16'b0000001100001000,
    16'b0000001101000011,
    16'b0000001000010000,
    16'b1111111110101000,
    16'b1111110011010100,
    16'b1111101010110101,
    16'b1111101001110010,
    16'b1111110011001101,
    16'b0000000111010011,
    16'b0000100011000111,
    16'b0001000001000000,
    16'b0001011010001010,
    16'b0001101000100001,
    16'b0001101000100001,
    16'b0001011010001010,
    16'b0001000001000000,
    16'b0000100011000111,
    16'b0000000111010011,
    16'b1111110011001101,
    16'b1111101001110010,
    16'b1111101010110101,
    16'b1111110011010100,
    16'b1111111110101000,
    16'b0000001000010000,
    16'b0000001101000011,
    16'b0000001100001000,
    16'b0000000110101111,
    16'b1111111111100100,
    16'b1111111001100010,
    16'b1111110110110010,
    16'b1111110111111011,
    16'b1111111100000100,
    16'b0000000001010001,
    16'b0000000101011010,
    16'b0000000111000001,
    16'b0000000101101110,
    16'b0000000010010100,
    16'b1111111110010101,
    16'b1111111011010110,
    16'b1111111010011110,
    16'b1111111011110101,
    16'b1111111110101110,
    16'b0000000001111001,
    16'b0000000100000011,
    16'b0000000100011101,
    16'b0000000011000101,
    16'b0000000000100101,
    16'b1111111110000010,
    16'b1111111100011100,
    16'b1111111100010111,
    16'b1111111101101111,
    16'b1111111111111011,
    16'b0000000010000001,
    16'b0000000011001101,
    16'b0000000011000100,
    16'b0000000001101110,
    16'b1111111111110001,
    16'b1111111110000000,
    16'b1111111101000111,
    16'b1111111101011010,
    16'b1111111110110000,
    16'b0000000000100110,
    16'b0000000010001110,
    16'b0000000011000010,
    16'b0000000010101111,
    16'b0000000001011111,
    16'b1111111111110000,
    16'b1111111110001101,
    16'b1111111101011101,
    16'b1111111101110111,
    16'b1111111111011000,
    16'b0000000001101001,
    16'b0000000100000101,
    16'b0000000110000110,
    16'b0000000111001110,
    16'b0000000111010010,
    16'b0000000110011000,
    16'b0000000100110010,
    16'b0000000010111011,
    16'b0000000001001101,
    16'b1111111111111000,
    16'b1111111111000110,
    16'b1111111110110011,
    16'b1111111110110111,
    16'b1111111111001000,
    16'b1111111111011101,
    16'b1111111111101110,
    16'b1111111111111001
};
